`ifndef INTER_F
`define INTER_F

interface inter_f(input logic clk, rst);
  
  bit data_in;
  logic full;
 
endinterface: inter_f
`endif