`ifndef MEM_AGENT_PKG
`define MEM_AGENT_PKG


package mem_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"



`include "sequence_item.sv"
`include "sequence.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"

endpackage
`endif
