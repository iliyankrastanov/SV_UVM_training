`ifndef MEM_TEST_LIST
`define MEM_TEST_LIST


package mem_test_list;

import uvm_pkg::*;
`include "uvm_macros.svh"

import mem_env_pkg::*;

`include "test.sv"

endpackage

`endif