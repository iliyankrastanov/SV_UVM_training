`ifndef MEM_ENV_PKG
`define MEM_ENV_PKG


package mem_env_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"


import mem_agent_pkg::*;

`include "environment.sv"

endpackage
`endif


